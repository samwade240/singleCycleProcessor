module programCounter_test();

reg clk,rst;
wire [7:0] count;


programCounter DUT(clk,rst,count);

initial
begin

	







end
endmodule
